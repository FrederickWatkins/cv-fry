import pipeline::*;
// Decoder
module idu (
    input decode_signals signals_in,

    output logic [4:0] rs1_addr,
    output logic [4:0] rs2_addr,
    output execute_signals signals_out
);
endmodule
