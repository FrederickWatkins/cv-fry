// Hazard controller